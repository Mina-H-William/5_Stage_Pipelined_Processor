LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY main IS
    GENERIC (

    );
    PORT (

    );
END main;

ARCHITECTURE Behavioral OF main IS

BEGIN
END Behavioral;