library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity main is
    generic (

    );
    Port (  
   
    );
end main;

architecture Behavioral of main is

begin


end Behavioral;


